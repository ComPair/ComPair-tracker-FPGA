../../vata_460p3/src/control_register_triggers.vhd